// Author:  Umberto Laghi
// Contact: umberto.laghi@studio.unibo.it
// Github:  @ubolakes

package trdb_pkg;
    // TODO: add correct length value
    localparam CAUSE_LEN = 5;
    localparam PRIV_LEN = 2; // depends on CPU implementation
    localparam INST_LEN = 32;
    localparam PTYPE_LEN = 4; // is it F + SF? spec not clear
    localparam P_LEN = 5;
    localparam PAYLOAD_LEN = 256;
    localparam TRIGGER_LEN = 4;
    localparam CTYPE_LEN = 2;
`ifdef TRDB_ARCH64 // 64bit arch specific parameters
    localparam XLEN = 64;
`else // 32bit arch
    localparam XLEN = 32;
`endif
    /* both archs parameters */
    // localparams for resync counter
    localparam CYCLE_MODE = 0;
    localparam PACKET_MODE = 1;
    // localparams for irreport and irdepth
    localparam CALL_COUNTER_SIZE = '0;
    localparam RETURN_STACK_SIZE = '0;
    // localparams for branch map - defined by spec
    localparam BRANCH_MAP_LEN = 31;
    localparam BRANCH_COUNT_LEN = 5;
    // localparams for filter mode
    localparam RANGE_MODE = 1'b0;
    localparam EQUAL_MODE = 1'b1;

// packet types
typedef enum logic[1:0] { 
    F_OPT_EXT       = 2'h0,
    F_DIFF_DELTA    = 2'h1,
    F_ADDR_ONLY     = 2'h2,
    F_SYNC          = 2'h3
} trdb_format_e;

// subformats available for type 3 packets (F_SYNC)
typedef enum logic[1:0] { 
    SF_START    = 2'h0,
    SF_TRAP     = 2'h1,
    SF_CONTEXT  = 2'h2,
    SF_SUPPORT  = 2'h3
} trdb_f_sync_subformat_e;

// subformats available for type 0 packets (F_OPT_EXT)
// used a struct for future extensions
typedef enum logic[0:0] {
    SF_PBC = 1'h0, // correctly predicted branches
    SF_JTC = 1'h1 // jump target cache in spec
} trdb_f_opt_ext_subformat_e;

// qual_status values necessary for format 3 subformat 3
// packet payload
typedef enum logic[1:0] {
    NO_CHANGE   = 2'h0,
    ENDED_REP   = 2'h1,
    TRACE_LOST  = 2'h2,
    ENDED_NTR   = 2'h3
} qual_status_e;

// enum that determines the ioptions values for
// format 3 subformat 3 packets
typedef enum logic[2:0] {
    DELTA_ADDRESS       = 3'h0,
    FULL_ADDRESS        = 3'h1,
    IMPLICIT_EXCEPTION  = 3'h2,
    SIJUMP              = 3'h3,
    IMPLICIT_RETURN     = 3'h4,
    BRANCH_PREDICTION   = 3'h5,
    JUMP_TARGET_CACHE   = 3'h6
} ioptions_e; // instruction trace options

// enum that expresses the packet format and 
// subformat to better readability
typedef enum logic[3:0] {
    F0SF0   = 4'h0,
    F0SF1   = 4'h1,
    F1      = 4'h4,
    F2      = 4'h8,
    F3SF0   = 4'hC,
    F3SF1   = 4'hD,
    F3SF2   = 4'hE,
    F3SF3   = 4'hF
} it_packet_type_e; // it stands for "instruction trace"

// defining packet structs for union
// format 3 subformat 0
typedef struct packed {
    trdb_f_sync_subformat_e subformat;
    logic                   branch;
    logic [PRIV_LEN-1:0]    priv_lvl;
    //logic [:0] time; // optional
    //logic [:0] context; // optional
    logic [XLEN-1:0]        address;
} f3_sf0_s;

// format 3 subformat 1
typedef struct packed {
    trdb_f_sync_subformat_e subformat;
    logic                   branch;
    logic [PRIV_LEN-1:0]    priv_lvl;
    //logic [:0] time; // optional
    //logic [:0] context; // optional
    logic [CAUSE_LEN-1:0]   ecause;
    logic                   interrupt;
    logic                   thaddr;
    logic [XLEN-1:0]        address;
    logic [XLEN-1:0]        tval;
} f3_sf1_s;

// format 3 subformat 2
typedef struct packed {
    trdb_f_sync_subformat_e subformat;
    logic [PRIV_LEN-1:0]    priv_lvl;
    //logic [:0] time; // optional
    //logic [:0] context; // optional
} f3_sf2_s;

// format 3 subformat 3
typedef struct packed {
    trdb_f_sync_subformat_e subformat;
    logic                   ienable;
    logic                   encoder_mode;
    qual_status_e           qual_status;
    ioptions_e              ioptions;
    //logic denable; // data trace support required
    //logic dloss; // data trace support required
    //logic [:0] doptions; // data trace support required
} f3_sf3_s;

// format 2
typedef struct packed {
    logic [XLEN-1:0]                address;
    logic                           notify;
    logic                           updiscon;
    logic                           irreport;
    logic [2**CALL_COUNTER_SIZE:0]  irdepth;
} f2_s;

// format 1 - branch_map w/address
typedef struct packed {
    logic [BRANCH_COUNT_LEN-1:0]    branches;
    logic [BRANCH_MAP_LEN-1:0]      branch_map;
    logic [XLEN-1:0]                address;
    logic                           notify;
    logic                           updiscon;
    logic                           irreport;
    logic [2**CALL_COUNTER_SIZE:0]  irdepth;
} f1_addr_s;

// format 1 - branch_map w/out address
typedef struct packed {
    logic [BRANCH_COUNT_LEN-1:0]    branches;
    logic [BRANCH_MAP_LEN-1:0]      branch_map;
} f1_no_addr_s;

// format 0 subformat 0 - branch_cnt w/out address
typedef struct packed {
    // TODO    
} f0_sf0_no_addr_s;

// format 0 subformat 0 - branch_cnt w/address
typedef struct packed {
    // TODO
} f0_sf0_addr_s;

// format 0 subformat 1 - jti w/branch_map
typedef struct packed {
    // TODO
} f0_sf1_map_s;

// format 0 subformat 1 - jti w/out branch_map
typedef struct packed {
    // TODO
} f0_sf1_no_map_s;

// payload union
typedef union packed {
    f3_sf0_s        f3_sf0;
    f3_sf1_s        f3_sf1;
    f3_sf2_s        f3_sf2;
    f3_sf3_s        f3_sf3;
    f2_s            f2;
    f1_addr_s       f1_addr;
    f1_no_addr_s    f1_no_addr;
    // TODO: add f0 packets
} packet_u;

// payload struct
typedef struct packed {
    trdb_format_e   format;
    packet_u        packet;
} packet_payload_s;

/*TODO:
    doptions struct for data tracing
    refer to page 36 of the spec */

/* Mask and match parameter for itype determination */
parameter MASK_BEQ = 32'h707f;
parameter MATCH_BEQ = 32'h63;
parameter MASK_BNE = 32'h707f;
parameter MATCH_BNE = 32'h1063;
parameter MASK_BLT = 32'h707f;
parameter MATCH_BLT = 32'h4063;
parameter MASK_BGE = 32'h707f;
parameter MATCH_BGE = 32'h5063;
parameter MASK_BLTU = 32'h707f;
parameter MATCH_BLTU = 32'h6063;
parameter MASK_BGEU = 32'h707f;
parameter MATCH_BGEU = 32'h7063;
parameter MASK_P_BNEIMM = 32'h707f;
parameter MATCH_P_BNEIMM = 32'h3063;
parameter MASK_P_BEQIMM = 32'h707f;
parameter MATCH_P_BEQIMM = 32'h2063;
parameter MASK_C_BEQZ = 32'he003;
parameter MATCH_C_BEQZ = 32'hc001;
parameter MASK_C_BNEZ = 32'he003;
parameter MATCH_C_BNEZ = 32'he001;
parameter MASK_C_JALR = 32'hf07f;
parameter MATCH_C_JALR = 32'h9002;
parameter MASK_RD = 32'hf80;
parameter MASK_C_JR = 32'hf07f;
parameter MATCH_C_JR = 32'h8002;
parameter MASK_JALR = 32'h707f;
parameter MATCH_JALR = 32'h67;
parameter MASK_MRET = 32'hffffffff;
parameter MATCH_MRET = 32'h30200073;
parameter MASK_SRET = 32'hffffffff;
parameter MATCH_SRET = 32'h10200073;
parameter MASK_URET = 32'hffffffff;
parameter MATCH_URET = 32'h200073;
parameter MASK_RS1 = 32'hf8000;
parameter MASK_IMM = 32'hfff00000;
parameter X_RA = 32'h1;
parameter OP_SH_RS1 = 32'd15;
parameter OP_SH_RD = 32'd7;




endpackage