/* PACKET EMITTER */
/*
it produces the packets for the output interface
*/

import trdb_pkg::*;

module trdb_packet_emitter
(
    // TO DO: add signals width

    input logic clk_i,
    input logic rst_ni,

    // necessary info to assemble packet
    input trdb_format_e packet_format_i,
    input trdb_subformat_e packet_subformat_i,

    // lc (last cycle) signals
    input logic lc_cause_i,
    input logic lc_tval,

    // tc (this cycle) signals
    input logic tc_cause_i,
    input logic tc_tval_i

    // nc (next cycle) signals


    // format 3 subformat 0 specific signals
    input logic is_branch_i,
    input logic is_branch_taken_i,
    input logic [PRIVLEN:0] priv_i,
    input logic [:0] time_i,    // optional
    input logic [:0] context_i, // optional
    input logic [XLEN-1:0] iaddr_i,

    // format 3 subformat 1 specific signals
    //input logic is_branch_i,
    //input logic is_branch_taken_i,
    //input logic [PRIVLEN:0] priv_i,
    //input logic [:0] time_i, // optional
    //input logic [:0] context_i, // optional
    input logic [CAUSELEN:0] ecause_i,
    input logic interrupt_i,
    input logic [XLEN-1:0] trap_handler_address_i, // is it the same as tvec?
    input logic [XLEN-1:0] epc_i,
    //input logic [XLEN-1:0]iaddr_i,
    input logic [TVALLEN:0] tval_i,

    // format 3 subformat 2 specific signals
    //input logic [PRIVLEN:0] priv_i,
    //input logic [:0] time_i, // optional
    //input logic [:0] context_i, // optional

    // format 3 subformat 3 specific signals
    input logic ienable_i, // trace encoder enabled
    input logic encoder_mode_i, // implementation specific, right now only branch trace supported (value==0). Hardwire to 0?
    //input logic [1:0] qual_status_i, // to be understood, generated by other signals?
    /*  it indicates the tracing has ended, it has two possible values: ended_rep and ended_ntr
        At page 37 of the specs there's a more accurate description*/
    // it doesn't require a dedicated input signal
    // because it's generated using other signals

    //input logic [:0] ioptions_i, // implementation specific
    // doesn't require an input, it must be created from other inputs
    /*  Run-time configuration bits for INSTRUCTION trace.
        Examples:
            - sequentially inferred jump: don't report the targets of sequentially inferable jumps
            - implicit return: don't report the targets of sequentially inferrable jumps
            - implicit exception: don't report function return addresses
            - branch prediction: branch predictor enabled (not supported in snitch)
            - jump target cache: enabled JTC (not supported in snitch)
            - full address: always output full addresses

        it requires info from the CSRs storing the values
    */
    //input logic seq_inferred_jump_i, // to implement
    input logic trace_implicit_ret_i,
    //input logic trace_implicit_exc_i, // to implement
    //input logic trace_branch_prediction_i, // not supported by snitch, hardwired to 0 (?)
    //input logic jump_target_cache_i, // not supported by snitch, hardwired to 0 (?)
    input logic trace_full_addr_i, // always output full address

    input logic denable_i, // DATA trace enabled, if supported
    // about DATA trace, in stand-by at the moment
    input logic dloss_i, // one or more DATA trace packets lost, if supported
    input logic [:0] doptions_i, // it's like ioptions, but for DATA trace


    // format 2 specific signals
    //input logic [XLEN-1:0] iaddr_i,
    /*  notify -> means the packet was requested by the cpu debug module
        not supported by snitch
        It requires an input from the priority module
    */ 
    input logic notify_i,
    /* updiscon ->  if it has a different value from notify,
                    means there was an exception/other flow 
                    changes during a loop.
                    This way the trace reconstruction is easier.
                    For a better description refer to page 38 of the spec
    */
    // most of the time these 2 values can be compressed
    //input logic lc_updiscon_i,

    input logic irreport_i,
    /*  the value of irreport is different from updiscon
        if this packet is reporting an instr that is the
        last one retired before an exception, interrupt, 
        priv change, resync.
        With this is also reported the traced nested calls, 
        that are counted if implicit_return mode is enabled
        (and available)
    */
    //input logic [:0] irdepth_i, // keeps count of the traced nested calls

    // format 1 specific signals
    /*  this format exists in two modes:
            - address, branch map
            - NO address, branch maps
        
        Their generation depends on the value of branches:
            - 0: no need for address
            - >0: address required
    */
    input logic [:0] branches_i, // in Robert implementation is called branch_cnt
    input logic [:0] branch_map_i, // in the packet it can change size to improve efficiency
    //input logic [XLEN-1:0] iaddr_i,
    //input logic notify_i,
    //input logic lc_updiscon_i,
    //input logic irreport_i, // same as format 2
    //input logic irdepth_i, // same as format 2
    

    // format 0 specific signals
    /*  This format can have two possible subformats:
            - subformat 0: number of correctly predicted branches
            - subformat 1: jump target cache index

    Since snitch does NOT support any of them,
    this format of packet is not necessary

    */
    //input logic [:0] branch_map_i,


    // outputs
    output logic [PTYPELEN:0]packet_type_o, // {packet_format, packet_subformat}
    output logic [PLEN:0] packet_length_o, // in bytes
    output logic [PAYLOADLEN:0] packet_payload_o,
    output logic packet_valid_o,

    /*outputs to perform reset resync counter
    and update/reset branch map.
    Question:   it should be done in this module or in
                the one choosing the packet format*/
    output logic branch_map_flush_o, // flushes the branch map
    output logic resync_timer_rst_o,  // not final
                                // understand how the Robert tracer does that

);
    
endmodule