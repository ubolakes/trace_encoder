/* PACKET EMITTER */
/*
it produces the packets for the output interface
*/

import trdb_pkg::*;

module trdb_packet_emitter
(
    input logic clk_i,
    input logic rst_ni,

    
);
    
endmodule