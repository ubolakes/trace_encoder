/* PACKET EMITTER */
/*
it produces the packets for the output interface
*/

import trdb_pkg::*;

module trdb_packet_emitter
(
    // TO DO: add signals width

    input logic clk_i,
    input logic rst_ni,

    input logic valid_i,

    // necessary info to assemble packet
    input trdb_format_e packet_format_i,
    input trdb_f_sync_subformat_e trdb_f_sync_subformat_i, // subformat for format 3
    //input trdb_f_opt_ext_subformat_e trdb_f_opt_ext_subformat_i, // non mandatory,subformat for format 0

    // lc (last cycle) signals
    input logic lc_cause_i,
    input logic lc_tval_i,

    // tc (this cycle) signals
    input logic tc_cause_i,
    input logic tc_tval_i,

    // nc (next cycle) signals


    // format 3 subformat 0 specific signals
    input logic is_branch_i,
    input logic is_branch_taken_i,
    input logic [PRIVLEN:0] priv_i,
    //input logic [:0] time_i,    // optional
    //input logic [:0] context_i, // optional
    input logic [XLEN-1:0] iaddr_i,
    input logic resync_timeout_i, // requested resync by the timer

    // format 3 subformat 1 specific signals
    //input logic is_branch_i,
    //input logic is_branch_taken_i,
    //input logic [PRIVLEN:0] priv_i,
    //input logic [:0] time_i, // optional
    //input logic [:0] context_i, // optional
    input logic cause_mux_i,
    /*  format 3 subformat 1 packets require sometimes lc_cause o tc_cause
        how do I discriminate them? Need another signal?
        The use of lc or tc values depends on a previous updiscon:
        combinatorial network that determines the ecause depending on
        the case.
        Idea:   output the ecause signal from trdb_priority, choosing
                between lc or tc*/
    input logic interrupt_i,
    input logic thaddr_i,
    input logic [XLEN-1:0] tvec_i, // trap handler address
    input logic [XLEN-1:0] epc_i,
    //input logic [XLEN-1:0]iaddr_i,
    input logic [TVALLEN:0] tval_i,

    // format 3 subformat 2 specific signals
    //input logic [PRIVLEN:0] priv_i,
    //input logic [:0] time_i, // optional
    //input logic [:0] context_i, // optional

    // format 3 subformat 3 specific signals
    input logic ienable_i, // trace encoder enabled
    input logic encoder_mode_i, // implementation specific, right now only branch trace supported (value==0). Hardwire to 0?
    input logic [1:0] qual_status_i, // to be understood, generated by other signals?
    /*  it indicates the tracing has ended, it has two possible values: ended_rep and ended_ntr
        At page 37 of the specs there's a more accurate description*/
    // it doesn't require a dedicated input signal
    // because it's generated using other signals

    input logic [:0] ioptions_i, // implementation specific
    /*  Run-time configuration bits for INSTRUCTION trace.
        These modes are optional, only the delta address is mandatory
        Examples:
            - sequentially inferred jump: don't report the targets of sequentially inferable jumps
            - implicit return: don't report the targets of sequentially inferrable jumps
            - implicit exception: don't report function return addresses
            - branch prediction: branch predictor enabled (not supported in snitch)
            - jump target cache: enabled JTC (not supported in snitch)
            - full address: always output full addresses

        it requires info from the CSRs storing the values
        For mandatory only modes it can be only 1
    */
    //input logic seq_inferred_jump_i, // to implement
    //input logic trace_implicit_ret_i, // implemented in Robert tracer
    //input logic trace_implicit_exc_i, // to implement
    //input logic trace_branch_prediction_i, // not supported by snitch, hardwired to 0 (?)
    //input logic jump_target_cache_i, // not supported by snitch, hardwired to 0 (?)
    //input logic trace_full_addr_i, // implemented in Robert tracer

    // about DATA trace, in stand-by at the moment
    //input logic denable_i, // DATA trace enabled, if supported
    //input logic dloss_i, // one or more DATA trace packets lost, if supported
    //input logic [:0] doptions_i, // it's like ioptions, but for DATA trace


    // format 2 specific signals
    //input logic [XLEN-1:0] iaddr_i,
    /*  notify -> means the packet was requested by the cpu trigger unit*/ 
    //input logic notify_i, // non mandatory
    
    /* updiscon ->  if it has a different value from notify,
                    means there was an exception/other flow 
                    changes during a loop.
                    This way the trace reconstruction is easier.
                    For a better description refer to page 38 of the spec
    */
    // most of the time these 2 values can be compressed
    input logic lc_updiscon_i,

    input logic irreport_i,
    /*  the value of irreport is different from updiscon
        if this packet is reporting an instr that is the
        last one retired before an exception, interrupt, 
        priv change, resync.
        With this is also reported the traced nested calls, 
        that are counted if implicit_return mode is enabled
        (and available)
    */
    //input logic [:0] irdepth_i, // keeps count of the traced nested calls

    // format 1 specific signals
    /*  this format exists in two modes:
            - address, branch map
            - NO address, branch maps
        
        Their generation depends on the value of branches:
            - 0: no need for address
            - >0: address required
    */
    input logic [:0] branches_i, // in Robert implementation is called branch_cnt
    input logic [:0] branch_map_i, // in the packet it can change size to improve efficiency
    //input logic [XLEN-1:0] iaddr_i,
    //input logic notify_i,
    //input logic lc_updiscon_i,
    //input logic irreport_i, // same as format 2
    //input logic irdepth_i, // same as format 2
    

    // format 0 specific signals
    /*  This format can have two possible subformats:
            - subformat 0: number of correctly predicted branches
            - subformat 1: jump target cache index

        Non mandatory, required support by the encoder.
    */
    //input logic [:0] branch_map_i,


    // outputs    ptypelen == 4?
    //output logic [PTYPELEN:0]packet_type_o, // {packet_format, packet_subformat}?
    //output logic [PLEN:0] payload_length_o, // in bytes
    /* this module produces only the packet payload
    that is the forwarded to the encapsulator that
    takes care of the type and length.*/
    output logic [PAYLOADLEN:0] packet_payload_o,
    output logic packet_valid_o, // asserted when a packet is generated

    output logic branch_map_flush_o, // branch map flushed after each request
    output logic resync_timer_rst_o,  // resets resync counter
);
    
    // internal signals
    logic branch;
    logic [XLEN-1:0] address;
    logic [CAUSELEN:0] ecause;
    logic [:0] diff_address;
    logic branch_map_flush_d, branch_map_flush_q;


    // assigning values
    assign branch = ~(is_branch_i && is_branch_taken_i);
    assign address = thaddr_i ? tvec_i : epc_i;
    assign ecause = cause_mux_i ? tc_cause_i : lc_cause_i;
    

    // combinatorial network to output packets
    always_comb begin : set_packet_bits
        // init values
        payload_length_o = '0; // in bytes, computed as the length in bit of (type+payload)/8
        packet_payload_o = '0;
        packet_valid_o = '0;
        
        if(valid_i) begin
            // flush the branch map
            /*  branch map flushing is done in the next cycle
                why? understand!*/
            branch_map_flush_d = '1;


            case(packet_format_i)

            F_SYNC: begin // format 3
                case(trdb_f_sync_subformat_i)

                SF_START: begin // subformat 0
                    packet_payload_o = {F_SYNC, F_START, branch, priv_i, /*time_i, context_i,*/ iaddr_i};
                    payload_length_o = (1 + PRIVLEN + /*TIMELEN: TBD + CONTEXTLEN: TBD*/ + XLEN-1)/8;
                    packet_valid_o = '1;
                end

                SF_TRAP: begin // subformat 1
                    packet_payload_o = {F_SYNC, SF_TRAP, branch, priv_i, /*time_i, context_i,*/ ecause, interrupt_i, thaddr_i, address, tval_i };
                    payload_length_o = ;
                    packet_valid_o = '1;
                end
                
                SF_CONTEXT: begin // subformat 2
                    packet_payload_o = {F_SYNC, SF_CONTEXT, priv_i/*,time_i, context_i*/};
                    payload_length_o = ;
                    packet_valid_o = '1;
                end
                
                SF_SUPPORT: begin // subformat 3
                    packet_payload_o = {F_SYNC, SF_SUPPORT, ienable_i, encoder_mode_i, qual_status_i, ioptions_i/*, denable_i, dloss_i, doptions_i*/};
                    payload_length_o = ;
                    packet_valid_o = '1;
                end
                endcase
            end


            F_ADDR_ONLY: begin // format 2
                packet_payload_o = {F_ADDR_ONLY, iaddr_i, /*notify_i,*/ lc_updiscon_i, irreport_i/*, irdepth_i*/};
                payload_length_o = ;
                packet_valid_o = '1;
            end


            F_DIFF_DELTA: begin // format 1
            /*  There can be two type of payloads for this format:
                1. address, branch map
                2. no address, branch map
                
                Type 1 payload is used when there has been at least
                one branch from last packet. This can be determined
                by the number of branches in the branch map.

                Type 2 payload is used when the address is not needed,
                for examples if the branch map is full.
            */
                if(branches_i < '31) begin // branch map not full - address
                    packet_payload_o = {F_DIFF_DELTA, branches_i, branch_map_i, iaddr_i, /*notify_i,*/ lc_updiscon_i, irreport_i/*, irdepth_i*/};
                    payload_length_o = ;
                end else /*if(branches_i == '31)*/ begin // branch map full - no address
                    packet_payload_o = {F_DIFF_DELTA, branches_i, branch_map_i};
                    payload_length_o = ;
                end
                packet_valid_o = '1;
            end


            F_OPT_EXT: begin // format 0
                /* requires non mandatory support for jtc and branch prediction
                case(trdb_f_opt_ext_subformat_i)
                SF_PBC: begin // subformat 0
                    packet_payload_o = {F_OPT_EXT, SF_PBC, etc..};
                    payload_length_o = ;
                    packet_valid_o = '1;
                end

                SF_JTC: begin // subformat 1
                    packet_payload_o = {F_OPT_EXT, SF_JTC, etc..};
                    payload_length_o = ;
                    packet_valid_o = '1;
                end
                endcase
                */
            end
            endcase
        
        end
    end


endmodule